// Project: SERICS - SANDSTORM
// Description: Set defines for CW305
// Author: Davide Bellizia <davide.bellizia@telsy.it>

`define CW305
`define ARTIX7
`define ARIANE_DATA_WIDTH 64

